** Profile: "rc_init_orcad_sch1-rc_init_bode"  [ u:\mes documents\mini projet 2015\travail_orcad\rc_init_orcad-pspicefiles\rc_init_orcad_sch1\rc_init_bode.sim ] 

** Creating circuit file "rc_init_bode.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\OrCAD\OrCAD_10.5\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 1000 10 1000k
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\rc_init_orcad_sch1.net" 


.END
